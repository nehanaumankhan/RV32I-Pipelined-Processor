`include "RISCV_PKG.vh"
module SCDP();
endmodule