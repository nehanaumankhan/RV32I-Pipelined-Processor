`include "RISCV_PKG.vh"
module alu_cu(
    input [6:0] opcode,
    input [2:0] funct3,
    input [6:0] funct7,
    output reg [3:0] alu_control
);

endmodule